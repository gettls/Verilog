module ex03(inX,inY,out);

    input inX,inY;
    output out;
    wire inX,inY;
    wire out;
    assign out = inX & inY;

endmodule