module ex02(in1, in2, in3, out1);

    input in1,in2,in3;
    output out1;

    wire in1,in2,in3;
    wire out1;

    assign out1=in1&in2&in3;
endmodule